VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO picorv32_woready
  CLASS BLOCK ;
  FOREIGN picorv32_woready ;
  ORIGIN 0.000 0.000 ;
  SIZE 586.335 BY 597.055 ;
  PIN VGND
    DIRECTION INPUT ;
    USE GROUND ;
    PORT
      LAYER met5 ;
        RECT 5.520 103.080 580.520 104.680 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 256.260 580.520 257.860 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 409.440 580.520 411.040 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 562.620 580.520 564.220 ;
    END
    PORT
      LAYER met4 ;
        RECT 97.840 10.640 99.440 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 251.440 10.640 253.040 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 405.040 10.640 406.640 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 558.640 10.640 560.240 585.040 ;
    END
  END VGND
  PIN VPWR
    DIRECTION INPUT ;
    USE POWER ;
    PORT
      LAYER met5 ;
        RECT 5.520 26.490 580.520 28.090 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 179.670 580.520 181.270 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 332.850 580.520 334.450 ;
    END
    PORT
      LAYER met5 ;
        RECT 5.520 486.030 580.520 487.630 ;
    END
    PORT
      LAYER met4 ;
        RECT 21.040 10.640 22.640 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 174.640 10.640 176.240 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 328.240 10.640 329.840 585.040 ;
    END
    PORT
      LAYER met4 ;
        RECT 481.840 10.640 483.440 585.040 ;
    END
  END VPWR
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 383.270 0.000 383.550 4.000 ;
    END
  END clk
  PIN eoi[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 12.970 593.055 13.250 597.055 ;
    END
  END eoi[0]
  PIN eoi[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 593.055 325.590 597.055 ;
    END
  END eoi[10]
  PIN eoi[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 593.055 100.190 597.055 ;
    END
  END eoi[11]
  PIN eoi[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 17.040 4.000 17.640 ;
    END
  END eoi[12]
  PIN eoi[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 309.440 586.335 310.040 ;
    END
  END eoi[13]
  PIN eoi[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 30.640 586.335 31.240 ;
    END
  END eoi[14]
  PIN eoi[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 267.350 593.055 267.630 597.055 ;
    END
  END eoi[15]
  PIN eoi[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 19.410 593.055 19.690 597.055 ;
    END
  END eoi[16]
  PIN eoi[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 196.510 0.000 196.790 4.000 ;
    END
  END eoi[17]
  PIN eoi[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 78.240 586.335 78.840 ;
    END
  END eoi[18]
  PIN eoi[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 523.640 586.335 524.240 ;
    END
  END eoi[19]
  PIN eoi[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 0.000 579.970 4.000 ;
    END
  END eoi[1]
  PIN eoi[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 57.840 4.000 58.440 ;
    END
  END eoi[20]
  PIN eoi[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 67.710 0.000 67.990 4.000 ;
    END
  END eoi[21]
  PIN eoi[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 71.440 586.335 72.040 ;
    END
  END eoi[22]
  PIN eoi[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 593.055 422.190 597.055 ;
    END
  END eoi[23]
  PIN eoi[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 106.350 0.000 106.630 4.000 ;
    END
  END eoi[24]
  PIN eoi[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 238.040 586.335 238.640 ;
    END
  END eoi[25]
  PIN eoi[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 183.640 4.000 184.240 ;
    END
  END eoi[26]
  PIN eoi[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 109.570 593.055 109.850 597.055 ;
    END
  END eoi[27]
  PIN eoi[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 180.240 586.335 180.840 ;
    END
  END eoi[28]
  PIN eoi[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 593.055 505.910 597.055 ;
    END
  END eoi[29]
  PIN eoi[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 479.870 0.000 480.150 4.000 ;
    END
  END eoi[2]
  PIN eoi[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 412.250 0.000 412.530 4.000 ;
    END
  END eoi[30]
  PIN eoi[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 64.640 4.000 65.240 ;
    END
  END eoi[31]
  PIN eoi[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 27.240 4.000 27.840 ;
    END
  END eoi[3]
  PIN eoi[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 495.970 0.000 496.250 4.000 ;
    END
  END eoi[4]
  PIN eoi[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 58.050 593.055 58.330 597.055 ;
    END
  END eoi[5]
  PIN eoi[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 363.840 586.335 364.440 ;
    END
  END eoi[6]
  PIN eoi[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 510.040 4.000 510.640 ;
    END
  END eoi[7]
  PIN eoi[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 431.570 593.055 431.850 597.055 ;
    END
  END eoi[8]
  PIN eoi[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 95.240 586.335 95.840 ;
    END
  END eoi[9]
  PIN irq[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 442.040 586.335 442.640 ;
    END
  END irq[0]
  PIN irq[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 0.000 534.890 4.000 ;
    END
  END irq[10]
  PIN irq[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 190.440 586.335 191.040 ;
    END
  END irq[11]
  PIN irq[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 570.030 0.000 570.310 4.000 ;
    END
  END irq[12]
  PIN irq[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 537.240 586.335 537.840 ;
    END
  END irq[13]
  PIN irq[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 156.440 586.335 157.040 ;
    END
  END irq[14]
  PIN irq[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 64.490 593.055 64.770 597.055 ;
    END
  END irq[15]
  PIN irq[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 593.055 332.030 597.055 ;
    END
  END irq[16]
  PIN irq[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 102.040 586.335 102.640 ;
    END
  END irq[17]
  PIN irq[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 582.910 593.055 583.190 597.055 ;
    END
  END irq[18]
  PIN irq[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 0.000 483.370 4.000 ;
    END
  END irq[19]
  PIN irq[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 595.040 4.000 595.640 ;
    END
  END irq[1]
  PIN irq[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 153.040 4.000 153.640 ;
    END
  END irq[20]
  PIN irq[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 540.640 4.000 541.240 ;
    END
  END irq[21]
  PIN irq[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 350.240 4.000 350.840 ;
    END
  END irq[22]
  PIN irq[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 146.240 4.000 146.840 ;
    END
  END irq[23]
  PIN irq[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 566.810 593.055 567.090 597.055 ;
    END
  END irq[24]
  PIN irq[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 340.040 4.000 340.640 ;
    END
  END irq[25]
  PIN irq[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 270.570 0.000 270.850 4.000 ;
    END
  END irq[26]
  PIN irq[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 561.040 586.335 561.640 ;
    END
  END irq[27]
  PIN irq[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 593.055 145.270 597.055 ;
    END
  END irq[28]
  PIN irq[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 64.640 586.335 65.240 ;
    END
  END irq[29]
  PIN irq[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 374.040 4.000 374.640 ;
    END
  END irq[2]
  PIN irq[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 285.640 4.000 286.240 ;
    END
  END irq[30]
  PIN irq[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 0.000 55.110 4.000 ;
    END
  END irq[31]
  PIN irq[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 593.055 116.290 597.055 ;
    END
  END irq[3]
  PIN irq[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 547.440 4.000 548.040 ;
    END
  END irq[4]
  PIN irq[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 421.640 4.000 422.240 ;
    END
  END irq[5]
  PIN irq[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 581.440 4.000 582.040 ;
    END
  END irq[6]
  PIN irq[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 593.055 138.830 597.055 ;
    END
  END irq[7]
  PIN irq[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 108.840 586.335 109.440 ;
    END
  END irq[8]
  PIN irq[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 265.240 4.000 265.840 ;
    END
  END irq[9]
  PIN mem_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 476.650 593.055 476.930 597.055 ;
    END
  END mem_addr[0]
  PIN mem_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 506.640 586.335 507.240 ;
    END
  END mem_addr[10]
  PIN mem_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 593.055 48.670 597.055 ;
    END
  END mem_addr[11]
  PIN mem_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 318.870 593.055 319.150 597.055 ;
    END
  END mem_addr[12]
  PIN mem_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 0.000 228.990 4.000 ;
    END
  END mem_addr[13]
  PIN mem_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 338.190 0.000 338.470 4.000 ;
    END
  END mem_addr[14]
  PIN mem_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 214.240 4.000 214.840 ;
    END
  END mem_addr[15]
  PIN mem_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 0.000 280.510 4.000 ;
    END
  END mem_addr[16]
  PIN mem_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 593.055 93.750 597.055 ;
    END
  END mem_addr[17]
  PIN mem_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 227.840 586.335 228.440 ;
    END
  END mem_addr[18]
  PIN mem_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 142.840 4.000 143.440 ;
    END
  END mem_addr[19]
  PIN mem_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 506.640 4.000 507.240 ;
    END
  END mem_addr[1]
  PIN mem_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 40.840 4.000 41.440 ;
    END
  END mem_addr[20]
  PIN mem_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 0.000 354.570 4.000 ;
    END
  END mem_addr[21]
  PIN mem_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 34.040 4.000 34.640 ;
    END
  END mem_addr[22]
  PIN mem_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 0.000 370.670 4.000 ;
    END
  END mem_addr[23]
  PIN mem_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 483.090 593.055 483.370 597.055 ;
    END
  END mem_addr[24]
  PIN mem_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 0.000 183.910 4.000 ;
    END
  END mem_addr[25]
  PIN mem_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 571.240 586.335 571.840 ;
    END
  END mem_addr[26]
  PIN mem_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 0.000 467.270 4.000 ;
    END
  END mem_addr[27]
  PIN mem_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 0.000 557.430 4.000 ;
    END
  END mem_addr[28]
  PIN mem_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 482.840 4.000 483.440 ;
    END
  END mem_addr[29]
  PIN mem_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 142.840 586.335 143.440 ;
    END
  END mem_addr[2]
  PIN mem_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 524.950 0.000 525.230 4.000 ;
    END
  END mem_addr[30]
  PIN mem_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 571.240 4.000 571.840 ;
    END
  END mem_addr[31]
  PIN mem_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 593.055 348.130 597.055 ;
    END
  END mem_addr[3]
  PIN mem_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 129.240 4.000 129.840 ;
    END
  END mem_addr[4]
  PIN mem_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 207.440 4.000 208.040 ;
    END
  END mem_addr[5]
  PIN mem_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 0.040 586.335 0.640 ;
    END
  END mem_addr[6]
  PIN mem_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 122.440 4.000 123.040 ;
    END
  END mem_addr[7]
  PIN mem_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 289.890 593.055 290.170 597.055 ;
    END
  END mem_addr[8]
  PIN mem_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 283.450 593.055 283.730 597.055 ;
    END
  END mem_addr[9]
  PIN mem_instr
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 312.430 593.055 312.710 597.055 ;
    END
  END mem_instr
  PIN mem_la_addr[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 323.040 586.335 323.640 ;
    END
  END mem_la_addr[0]
  PIN mem_la_addr[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 593.055 3.590 597.055 ;
    END
  END mem_la_addr[10]
  PIN mem_la_addr[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 199.730 593.055 200.010 597.055 ;
    END
  END mem_la_addr[11]
  PIN mem_la_addr[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 296.330 593.055 296.610 597.055 ;
    END
  END mem_la_addr[12]
  PIN mem_la_addr[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 593.055 303.050 597.055 ;
    END
  END mem_la_addr[13]
  PIN mem_la_addr[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 593.055 377.110 597.055 ;
    END
  END mem_la_addr[14]
  PIN mem_la_addr[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 238.040 4.000 238.640 ;
    END
  END mem_la_addr[15]
  PIN mem_la_addr[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 138.550 0.000 138.830 4.000 ;
    END
  END mem_la_addr[16]
  PIN mem_la_addr[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 367.240 4.000 367.840 ;
    END
  END mem_la_addr[17]
  PIN mem_la_addr[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 554.240 4.000 554.840 ;
    END
  END mem_la_addr[18]
  PIN mem_la_addr[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 0.000 206.450 4.000 ;
    END
  END mem_la_addr[19]
  PIN mem_la_addr[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 0.000 167.810 4.000 ;
    END
  END mem_la_addr[1]
  PIN mem_la_addr[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 593.055 257.970 597.055 ;
    END
  END mem_la_addr[20]
  PIN mem_la_addr[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 333.240 4.000 333.840 ;
    END
  END mem_la_addr[21]
  PIN mem_la_addr[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 341.410 593.055 341.690 597.055 ;
    END
  END mem_la_addr[22]
  PIN mem_la_addr[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 80.590 593.055 80.870 597.055 ;
    END
  END mem_la_addr[23]
  PIN mem_la_addr[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 521.730 593.055 522.010 597.055 ;
    END
  END mem_la_addr[24]
  PIN mem_la_addr[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 377.440 586.335 378.040 ;
    END
  END mem_la_addr[25]
  PIN mem_la_addr[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 523.640 4.000 524.240 ;
    END
  END mem_la_addr[26]
  PIN mem_la_addr[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 35.510 593.055 35.790 597.055 ;
    END
  END mem_la_addr[27]
  PIN mem_la_addr[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 85.040 586.335 85.640 ;
    END
  END mem_la_addr[28]
  PIN mem_la_addr[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 214.240 586.335 214.840 ;
    END
  END mem_la_addr[29]
  PIN mem_la_addr[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 231.240 586.335 231.840 ;
    END
  END mem_la_addr[2]
  PIN mem_la_addr[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 593.055 393.210 597.055 ;
    END
  END mem_la_addr[30]
  PIN mem_la_addr[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 593.055 489.810 597.055 ;
    END
  END mem_la_addr[31]
  PIN mem_la_addr[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 6.530 593.055 6.810 597.055 ;
    END
  END mem_la_addr[3]
  PIN mem_la_addr[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 447.670 593.055 447.950 597.055 ;
    END
  END mem_la_addr[4]
  PIN mem_la_addr[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 489.640 586.335 490.240 ;
    END
  END mem_la_addr[5]
  PIN mem_la_addr[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 173.970 0.000 174.250 4.000 ;
    END
  END mem_la_addr[6]
  PIN mem_la_addr[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 112.240 586.335 112.840 ;
    END
  END mem_la_addr[7]
  PIN mem_la_addr[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 469.240 4.000 469.840 ;
    END
  END mem_la_addr[8]
  PIN mem_la_addr[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 132.640 586.335 133.240 ;
    END
  END mem_la_addr[9]
  PIN mem_la_read
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 515.290 593.055 515.570 597.055 ;
    END
  END mem_la_read
  PIN mem_la_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 425.040 586.335 425.640 ;
    END
  END mem_la_wdata[0]
  PIN mem_la_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 414.840 4.000 415.440 ;
    END
  END mem_la_wdata[10]
  PIN mem_la_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 103.130 593.055 103.410 597.055 ;
    END
  END mem_la_wdata[11]
  PIN mem_la_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 421.910 0.000 422.190 4.000 ;
    END
  END mem_la_wdata[12]
  PIN mem_la_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 392.930 0.000 393.210 4.000 ;
    END
  END mem_la_wdata[13]
  PIN mem_la_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 228.710 593.055 228.990 597.055 ;
    END
  END mem_la_wdata[14]
  PIN mem_la_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 248.030 0.000 248.310 4.000 ;
    END
  END mem_la_wdata[15]
  PIN mem_la_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 537.830 593.055 538.110 597.055 ;
    END
  END mem_la_wdata[16]
  PIN mem_la_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 593.055 274.070 597.055 ;
    END
  END mem_la_wdata[17]
  PIN mem_la_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 0.000 190.350 4.000 ;
    END
  END mem_la_wdata[18]
  PIN mem_la_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 264.130 0.000 264.410 4.000 ;
    END
  END mem_la_wdata[19]
  PIN mem_la_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 418.240 586.335 418.840 ;
    END
  END mem_la_wdata[1]
  PIN mem_la_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 241.440 4.000 242.040 ;
    END
  END mem_la_wdata[20]
  PIN mem_la_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 302.640 4.000 303.240 ;
    END
  END mem_la_wdata[21]
  PIN mem_la_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 411.440 586.335 412.040 ;
    END
  END mem_la_wdata[22]
  PIN mem_la_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 316.240 4.000 316.840 ;
    END
  END mem_la_wdata[23]
  PIN mem_la_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 344.630 0.000 344.910 4.000 ;
    END
  END mem_la_wdata[24]
  PIN mem_la_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 462.440 4.000 463.040 ;
    END
  END mem_la_wdata[25]
  PIN mem_la_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 112.240 4.000 112.840 ;
    END
  END mem_la_wdata[26]
  PIN mem_la_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 135.330 0.000 135.610 4.000 ;
    END
  END mem_la_wdata[27]
  PIN mem_la_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 593.055 251.530 597.055 ;
    END
  END mem_la_wdata[28]
  PIN mem_la_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 257.690 0.000 257.970 4.000 ;
    END
  END mem_la_wdata[29]
  PIN mem_la_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 278.840 4.000 279.440 ;
    END
  END mem_la_wdata[2]
  PIN mem_la_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 593.055 77.650 597.055 ;
    END
  END mem_la_wdata[30]
  PIN mem_la_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 136.040 586.335 136.640 ;
    END
  END mem_la_wdata[31]
  PIN mem_la_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 166.640 4.000 167.240 ;
    END
  END mem_la_wdata[3]
  PIN mem_la_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 376.830 0.000 377.110 4.000 ;
    END
  END mem_la_wdata[4]
  PIN mem_la_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 578.040 586.335 578.640 ;
    END
  END mem_la_wdata[5]
  PIN mem_la_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 202.950 0.000 203.230 4.000 ;
    END
  END mem_la_wdata[6]
  PIN mem_la_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 411.440 4.000 412.040 ;
    END
  END mem_la_wdata[7]
  PIN mem_la_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 261.840 4.000 262.440 ;
    END
  END mem_la_wdata[8]
  PIN mem_la_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 486.240 4.000 486.840 ;
    END
  END mem_la_wdata[9]
  PIN mem_la_write
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 593.055 460.830 597.055 ;
    END
  END mem_la_write
  PIN mem_la_wstrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 533.840 4.000 534.440 ;
    END
  END mem_la_wstrb[0]
  PIN mem_la_wstrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 261.840 586.335 262.440 ;
    END
  END mem_la_wstrb[1]
  PIN mem_la_wstrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 154.650 593.055 154.930 597.055 ;
    END
  END mem_la_wstrb[2]
  PIN mem_la_wstrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 319.640 4.000 320.240 ;
    END
  END mem_la_wstrb[3]
  PIN mem_rdata[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 496.440 586.335 497.040 ;
    END
  END mem_rdata[0]
  PIN mem_rdata[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 260.910 593.055 261.190 597.055 ;
    END
  END mem_rdata[10]
  PIN mem_rdata[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 278.840 586.335 279.440 ;
    END
  END mem_rdata[11]
  PIN mem_rdata[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 354.290 593.055 354.570 597.055 ;
    END
  END mem_rdata[12]
  PIN mem_rdata[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 405.810 0.000 406.090 4.000 ;
    END
  END mem_rdata[13]
  PIN mem_rdata[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 445.440 4.000 446.040 ;
    END
  END mem_rdata[14]
  PIN mem_rdata[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 183.630 593.055 183.910 597.055 ;
    END
  END mem_rdata[15]
  PIN mem_rdata[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 221.040 586.335 221.640 ;
    END
  END mem_rdata[16]
  PIN mem_rdata[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 544.040 586.335 544.640 ;
    END
  END mem_rdata[17]
  PIN mem_rdata[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 380.840 4.000 381.440 ;
    END
  END mem_rdata[18]
  PIN mem_rdata[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 119.040 4.000 119.640 ;
    END
  END mem_rdata[19]
  PIN mem_rdata[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 272.040 4.000 272.640 ;
    END
  END mem_rdata[1]
  PIN mem_rdata[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 299.550 0.000 299.830 4.000 ;
    END
  END mem_rdata[20]
  PIN mem_rdata[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 255.040 586.335 255.640 ;
    END
  END mem_rdata[21]
  PIN mem_rdata[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 584.840 586.335 585.440 ;
    END
  END mem_rdata[22]
  PIN mem_rdata[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 401.240 586.335 401.840 ;
    END
  END mem_rdata[23]
  PIN mem_rdata[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 346.840 586.335 347.440 ;
    END
  END mem_rdata[24]
  PIN mem_rdata[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 0.000 161.370 4.000 ;
    END
  END mem_rdata[25]
  PIN mem_rdata[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 593.055 438.290 597.055 ;
    END
  END mem_rdata[26]
  PIN mem_rdata[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 302.770 0.000 303.050 4.000 ;
    END
  END mem_rdata[27]
  PIN mem_rdata[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 222.270 593.055 222.550 597.055 ;
    END
  END mem_rdata[28]
  PIN mem_rdata[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 77.370 0.000 77.650 4.000 ;
    END
  END mem_rdata[29]
  PIN mem_rdata[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 452.240 586.335 452.840 ;
    END
  END mem_rdata[2]
  PIN mem_rdata[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 241.590 0.000 241.870 4.000 ;
    END
  END mem_rdata[30]
  PIN mem_rdata[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 71.440 4.000 72.040 ;
    END
  END mem_rdata[31]
  PIN mem_rdata[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 248.240 4.000 248.840 ;
    END
  END mem_rdata[3]
  PIN mem_rdata[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 215.830 593.055 216.110 597.055 ;
    END
  END mem_rdata[4]
  PIN mem_rdata[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 363.950 593.055 364.230 597.055 ;
    END
  END mem_rdata[5]
  PIN mem_rdata[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 593.055 32.570 597.055 ;
    END
  END mem_rdata[6]
  PIN mem_rdata[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 273.790 0.000 274.070 4.000 ;
    END
  END mem_rdata[7]
  PIN mem_rdata[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 334.970 593.055 335.250 597.055 ;
    END
  END mem_rdata[8]
  PIN mem_rdata[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 81.640 4.000 82.240 ;
    END
  END mem_rdata[9]
  PIN mem_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 207.440 586.335 208.040 ;
    END
  END mem_valid
  PIN mem_wdata[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 435.240 4.000 435.840 ;
    END
  END mem_wdata[0]
  PIN mem_wdata[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 193.840 4.000 194.440 ;
    END
  END mem_wdata[10]
  PIN mem_wdata[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 176.840 4.000 177.440 ;
    END
  END mem_wdata[11]
  PIN mem_wdata[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 547.490 0.000 547.770 4.000 ;
    END
  END mem_wdata[12]
  PIN mem_wdata[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 95.240 4.000 95.840 ;
    END
  END mem_wdata[13]
  PIN mem_wdata[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 482.840 586.335 483.440 ;
    END
  END mem_wdata[14]
  PIN mem_wdata[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 32.290 0.000 32.570 4.000 ;
    END
  END mem_wdata[15]
  PIN mem_wdata[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 0.000 235.430 4.000 ;
    END
  END mem_wdata[16]
  PIN mem_wdata[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 387.640 4.000 388.240 ;
    END
  END mem_wdata[17]
  PIN mem_wdata[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 518.510 0.000 518.790 4.000 ;
    END
  END mem_wdata[18]
  PIN mem_wdata[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 438.640 4.000 439.240 ;
    END
  END mem_wdata[19]
  PIN mem_wdata[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 370.390 593.055 370.670 597.055 ;
    END
  END mem_wdata[1]
  PIN mem_wdata[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 0.000 512.350 4.000 ;
    END
  END mem_wdata[20]
  PIN mem_wdata[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 404.640 4.000 405.240 ;
    END
  END mem_wdata[21]
  PIN mem_wdata[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 47.640 586.335 48.240 ;
    END
  END mem_wdata[22]
  PIN mem_wdata[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 224.440 4.000 225.040 ;
    END
  END mem_wdata[23]
  PIN mem_wdata[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 231.240 4.000 231.840 ;
    END
  END mem_wdata[24]
  PIN mem_wdata[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 315.650 0.000 315.930 4.000 ;
    END
  END mem_wdata[25]
  PIN mem_wdata[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 357.040 4.000 357.640 ;
    END
  END mem_wdata[26]
  PIN mem_wdata[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 238.370 593.055 238.650 597.055 ;
    END
  END mem_wdata[27]
  PIN mem_wdata[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 119.040 586.335 119.640 ;
    END
  END mem_wdata[28]
  PIN mem_wdata[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 217.640 4.000 218.240 ;
    END
  END mem_wdata[29]
  PIN mem_wdata[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 578.040 4.000 578.640 ;
    END
  END mem_wdata[2]
  PIN mem_wdata[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 520.240 586.335 520.840 ;
    END
  END mem_wdata[30]
  PIN mem_wdata[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 493.040 4.000 493.640 ;
    END
  END mem_wdata[31]
  PIN mem_wdata[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 309.440 4.000 310.040 ;
    END
  END mem_wdata[3]
  PIN mem_wdata[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 151.430 0.000 151.710 4.000 ;
    END
  END mem_wdata[4]
  PIN mem_wdata[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 489.530 0.000 489.810 4.000 ;
    END
  END mem_wdata[5]
  PIN mem_wdata[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 23.840 586.335 24.440 ;
    END
  END mem_wdata[6]
  PIN mem_wdata[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 428.440 4.000 429.040 ;
    END
  END mem_wdata[7]
  PIN mem_wdata[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 579.690 593.055 579.970 597.055 ;
    END
  END mem_wdata[8]
  PIN mem_wdata[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 360.730 0.000 361.010 4.000 ;
    END
  END mem_wdata[9]
  PIN mem_wstrb[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 268.640 586.335 269.240 ;
    END
  END mem_wstrb[0]
  PIN mem_wstrb[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 204.040 586.335 204.640 ;
    END
  END mem_wstrb[1]
  PIN mem_wstrb[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 404.640 586.335 405.240 ;
    END
  END mem_wstrb[2]
  PIN mem_wstrb[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 316.240 586.335 316.840 ;
    END
  END mem_wstrb[3]
  PIN pcpi_insn[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 244.810 593.055 245.090 597.055 ;
    END
  END pcpi_insn[0]
  PIN pcpi_insn[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 329.840 586.335 330.440 ;
    END
  END pcpi_insn[10]
  PIN pcpi_insn[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 23.840 4.000 24.440 ;
    END
  END pcpi_insn[11]
  PIN pcpi_insn[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 502.410 0.000 502.690 4.000 ;
    END
  END pcpi_insn[12]
  PIN pcpi_insn[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 83.810 0.000 84.090 4.000 ;
    END
  END pcpi_insn[13]
  PIN pcpi_insn[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 74.840 4.000 75.440 ;
    END
  END pcpi_insn[14]
  PIN pcpi_insn[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 450.890 0.000 451.170 4.000 ;
    END
  END pcpi_insn[15]
  PIN pcpi_insn[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 37.440 586.335 38.040 ;
    END
  END pcpi_insn[16]
  PIN pcpi_insn[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 132.110 593.055 132.390 597.055 ;
    END
  END pcpi_insn[17]
  PIN pcpi_insn[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 557.150 593.055 557.430 597.055 ;
    END
  END pcpi_insn[18]
  PIN pcpi_insn[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 593.055 122.730 597.055 ;
    END
  END pcpi_insn[19]
  PIN pcpi_insn[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 459.040 4.000 459.640 ;
    END
  END pcpi_insn[1]
  PIN pcpi_insn[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 157.870 0.000 158.150 4.000 ;
    END
  END pcpi_insn[20]
  PIN pcpi_insn[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 564.440 4.000 565.040 ;
    END
  END pcpi_insn[21]
  PIN pcpi_insn[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 505.630 0.000 505.910 4.000 ;
    END
  END pcpi_insn[22]
  PIN pcpi_insn[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 593.055 415.750 597.055 ;
    END
  END pcpi_insn[23]
  PIN pcpi_insn[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 99.910 0.000 100.190 4.000 ;
    END
  END pcpi_insn[24]
  PIN pcpi_insn[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 299.240 586.335 299.840 ;
    END
  END pcpi_insn[25]
  PIN pcpi_insn[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 554.240 586.335 554.840 ;
    END
  END pcpi_insn[26]
  PIN pcpi_insn[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 591.640 586.335 592.240 ;
    END
  END pcpi_insn[27]
  PIN pcpi_insn[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 499.840 586.335 500.440 ;
    END
  END pcpi_insn[28]
  PIN pcpi_insn[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 476.040 586.335 476.640 ;
    END
  END pcpi_insn[29]
  PIN pcpi_insn[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 472.640 586.335 473.240 ;
    END
  END pcpi_insn[2]
  PIN pcpi_insn[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 255.040 4.000 255.640 ;
    END
  END pcpi_insn[30]
  PIN pcpi_insn[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 534.610 593.055 534.890 597.055 ;
    END
  END pcpi_insn[31]
  PIN pcpi_insn[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 16.190 0.000 16.470 4.000 ;
    END
  END pcpi_insn[3]
  PIN pcpi_insn[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 3.310 0.000 3.590 4.000 ;
    END
  END pcpi_insn[4]
  PIN pcpi_insn[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 593.055 26.130 597.055 ;
    END
  END pcpi_insn[5]
  PIN pcpi_insn[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 293.110 0.000 293.390 4.000 ;
    END
  END pcpi_insn[6]
  PIN pcpi_insn[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 6.840 586.335 7.440 ;
    END
  END pcpi_insn[7]
  PIN pcpi_insn[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 573.250 593.055 573.530 597.055 ;
    END
  END pcpi_insn[8]
  PIN pcpi_insn[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 54.440 586.335 55.040 ;
    END
  END pcpi_insn[9]
  PIN pcpi_rd[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 235.150 593.055 235.430 597.055 ;
    END
  END pcpi_rd[0]
  PIN pcpi_rd[10]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 391.040 4.000 391.640 ;
    END
  END pcpi_rd[10]
  PIN pcpi_rd[11]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 112.790 0.000 113.070 4.000 ;
    END
  END pcpi_rd[11]
  PIN pcpi_rd[12]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 251.250 0.000 251.530 4.000 ;
    END
  END pcpi_rd[12]
  PIN pcpi_rd[13]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 499.190 593.055 499.470 597.055 ;
    END
  END pcpi_rd[13]
  PIN pcpi_rd[14]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 159.840 4.000 160.440 ;
    END
  END pcpi_rd[14]
  PIN pcpi_rd[15]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 0.000 212.890 4.000 ;
    END
  END pcpi_rd[15]
  PIN pcpi_rd[16]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 452.240 4.000 452.840 ;
    END
  END pcpi_rd[16]
  PIN pcpi_rd[17]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 275.440 586.335 276.040 ;
    END
  END pcpi_rd[17]
  PIN pcpi_rd[18]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 387.640 586.335 388.240 ;
    END
  END pcpi_rd[18]
  PIN pcpi_rd[19]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 438.010 0.000 438.290 4.000 ;
    END
  END pcpi_rd[19]
  PIN pcpi_rd[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 206.170 593.055 206.450 597.055 ;
    END
  END pcpi_rd[1]
  PIN pcpi_rd[20]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 563.590 0.000 563.870 4.000 ;
    END
  END pcpi_rd[20]
  PIN pcpi_rd[21]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 370.640 586.335 371.240 ;
    END
  END pcpi_rd[21]
  PIN pcpi_rd[22]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 98.640 4.000 99.240 ;
    END
  END pcpi_rd[22]
  PIN pcpi_rd[23]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 292.440 586.335 293.040 ;
    END
  END pcpi_rd[23]
  PIN pcpi_rd[24]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 434.790 0.000 435.070 4.000 ;
    END
  END pcpi_rd[24]
  PIN pcpi_rd[25]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 593.055 528.450 597.055 ;
    END
  END pcpi_rd[25]
  PIN pcpi_rd[26]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 40.840 586.335 41.440 ;
    END
  END pcpi_rd[26]
  PIN pcpi_rd[27]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 357.510 593.055 357.790 597.055 ;
    END
  END pcpi_rd[27]
  PIN pcpi_rd[28]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 528.170 0.000 528.450 4.000 ;
    END
  END pcpi_rd[28]
  PIN pcpi_rd[29]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 161.090 593.055 161.370 597.055 ;
    END
  END pcpi_rd[29]
  PIN pcpi_rd[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 0.000 71.210 4.000 ;
    END
  END pcpi_rd[2]
  PIN pcpi_rd[30]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 3.440 4.000 4.040 ;
    END
  END pcpi_rd[30]
  PIN pcpi_rd[31]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 588.240 4.000 588.840 ;
    END
  END pcpi_rd[31]
  PIN pcpi_rd[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 380.840 586.335 381.440 ;
    END
  END pcpi_rd[3]
  PIN pcpi_rd[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 144.990 0.000 145.270 4.000 ;
    END
  END pcpi_rd[4]
  PIN pcpi_rd[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 541.050 0.000 541.330 4.000 ;
    END
  END pcpi_rd[5]
  PIN pcpi_rd[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 190.070 593.055 190.350 597.055 ;
    END
  END pcpi_rd[6]
  PIN pcpi_rd[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 512.070 593.055 512.350 597.055 ;
    END
  END pcpi_rd[7]
  PIN pcpi_rd[8]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 448.840 586.335 449.440 ;
    END
  END pcpi_rd[8]
  PIN pcpi_rd[9]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 167.530 593.055 167.810 597.055 ;
    END
  END pcpi_rd[9]
  PIN pcpi_ready
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 88.440 4.000 89.040 ;
    END
  END pcpi_ready
  PIN pcpi_rs1[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 88.440 586.335 89.040 ;
    END
  END pcpi_rs1[0]
  PIN pcpi_rs1[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 125.670 593.055 125.950 597.055 ;
    END
  END pcpi_rs1[10]
  PIN pcpi_rs1[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 197.240 586.335 197.840 ;
    END
  END pcpi_rs1[11]
  PIN pcpi_rs1[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 593.055 399.650 597.055 ;
    END
  END pcpi_rs1[12]
  PIN pcpi_rs1[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 280.230 593.055 280.510 597.055 ;
    END
  END pcpi_rs1[13]
  PIN pcpi_rs1[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 54.830 593.055 55.110 597.055 ;
    END
  END pcpi_rs1[14]
  PIN pcpi_rs1[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 48.390 0.000 48.670 4.000 ;
    END
  END pcpi_rs1[15]
  PIN pcpi_rs1[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 322.090 0.000 322.370 4.000 ;
    END
  END pcpi_rs1[16]
  PIN pcpi_rs1[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 428.440 586.335 429.040 ;
    END
  END pcpi_rs1[17]
  PIN pcpi_rs1[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 394.440 586.335 395.040 ;
    END
  END pcpi_rs1[18]
  PIN pcpi_rs1[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 367.170 0.000 367.450 4.000 ;
    END
  END pcpi_rs1[19]
  PIN pcpi_rs1[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 343.440 4.000 344.040 ;
    END
  END pcpi_rs1[1]
  PIN pcpi_rs1[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 173.440 586.335 174.040 ;
    END
  END pcpi_rs1[20]
  PIN pcpi_rs1[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 0.000 550.990 4.000 ;
    END
  END pcpi_rs1[21]
  PIN pcpi_rs1[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 47.640 4.000 48.240 ;
    END
  END pcpi_rs1[22]
  PIN pcpi_rs1[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 550.710 593.055 550.990 597.055 ;
    END
  END pcpi_rs1[23]
  PIN pcpi_rs1[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 325.310 0.000 325.590 4.000 ;
    END
  END pcpi_rs1[24]
  PIN pcpi_rs1[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 460.550 0.000 460.830 4.000 ;
    END
  END pcpi_rs1[25]
  PIN pcpi_rs1[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 125.840 586.335 126.440 ;
    END
  END pcpi_rs1[26]
  PIN pcpi_rs1[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 87.030 593.055 87.310 597.055 ;
    END
  END pcpi_rs1[27]
  PIN pcpi_rs1[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 105.440 4.000 106.040 ;
    END
  END pcpi_rs1[28]
  PIN pcpi_rs1[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 61.270 0.000 61.550 4.000 ;
    END
  END pcpi_rs1[29]
  PIN pcpi_rs1[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 212.610 593.055 212.890 597.055 ;
    END
  END pcpi_rs1[2]
  PIN pcpi_rs1[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 340.040 586.335 340.640 ;
    END
  END pcpi_rs1[30]
  PIN pcpi_rs1[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 567.840 586.335 568.440 ;
    END
  END pcpi_rs1[31]
  PIN pcpi_rs1[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 225.490 0.000 225.770 4.000 ;
    END
  END pcpi_rs1[3]
  PIN pcpi_rs1[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 470.210 593.055 470.490 597.055 ;
    END
  END pcpi_rs1[4]
  PIN pcpi_rs1[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 244.840 586.335 245.440 ;
    END
  END pcpi_rs1[5]
  PIN pcpi_rs1[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 0.000 444.730 4.000 ;
    END
  END pcpi_rs1[6]
  PIN pcpi_rs1[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 454.110 593.055 454.390 597.055 ;
    END
  END pcpi_rs1[7]
  PIN pcpi_rs1[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 428.350 0.000 428.630 4.000 ;
    END
  END pcpi_rs1[8]
  PIN pcpi_rs1[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 295.840 4.000 296.440 ;
    END
  END pcpi_rs1[9]
  PIN pcpi_rs2[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 25.850 0.000 26.130 4.000 ;
    END
  END pcpi_rs2[0]
  PIN pcpi_rs2[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 576.470 0.000 576.750 4.000 ;
    END
  END pcpi_rs2[10]
  PIN pcpi_rs2[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 149.640 586.335 150.240 ;
    END
  END pcpi_rs2[11]
  PIN pcpi_rs2[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 193.290 593.055 193.570 597.055 ;
    END
  END pcpi_rs2[12]
  PIN pcpi_rs2[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 513.440 586.335 514.040 ;
    END
  END pcpi_rs2[13]
  PIN pcpi_rs2[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 476.040 4.000 476.640 ;
    END
  END pcpi_rs2[14]
  PIN pcpi_rs2[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 516.840 4.000 517.440 ;
    END
  END pcpi_rs2[15]
  PIN pcpi_rs2[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 10.240 4.000 10.840 ;
    END
  END pcpi_rs2[16]
  PIN pcpi_rs2[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 22.630 0.000 22.910 4.000 ;
    END
  END pcpi_rs2[17]
  PIN pcpi_rs2[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 122.450 0.000 122.730 4.000 ;
    END
  END pcpi_rs2[18]
  PIN pcpi_rs2[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 306.040 586.335 306.640 ;
    END
  END pcpi_rs2[19]
  PIN pcpi_rs2[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 331.750 0.000 332.030 4.000 ;
    END
  END pcpi_rs2[1]
  PIN pcpi_rs2[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 402.590 593.055 402.870 597.055 ;
    END
  END pcpi_rs2[20]
  PIN pcpi_rs2[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 544.270 593.055 544.550 597.055 ;
    END
  END pcpi_rs2[21]
  PIN pcpi_rs2[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 41.950 593.055 42.230 597.055 ;
    END
  END pcpi_rs2[22]
  PIN pcpi_rs2[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 90.250 0.000 90.530 4.000 ;
    END
  END pcpi_rs2[23]
  PIN pcpi_rs2[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 353.640 586.335 354.240 ;
    END
  END pcpi_rs2[24]
  PIN pcpi_rs2[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 560.370 593.055 560.650 597.055 ;
    END
  END pcpi_rs2[25]
  PIN pcpi_rs2[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 363.840 4.000 364.440 ;
    END
  END pcpi_rs2[26]
  PIN pcpi_rs2[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 465.840 586.335 466.440 ;
    END
  END pcpi_rs2[27]
  PIN pcpi_rs2[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 183.640 586.335 184.240 ;
    END
  END pcpi_rs2[28]
  PIN pcpi_rs2[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 399.370 0.000 399.650 4.000 ;
    END
  END pcpi_rs2[29]
  PIN pcpi_rs2[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 492.750 593.055 493.030 597.055 ;
    END
  END pcpi_rs2[2]
  PIN pcpi_rs2[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 148.210 593.055 148.490 597.055 ;
    END
  END pcpi_rs2[30]
  PIN pcpi_rs2[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 180.410 0.000 180.690 4.000 ;
    END
  END pcpi_rs2[31]
  PIN pcpi_rs2[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 357.040 586.335 357.640 ;
    END
  END pcpi_rs2[3]
  PIN pcpi_rs2[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 473.430 0.000 473.710 4.000 ;
    END
  END pcpi_rs2[4]
  PIN pcpi_rs2[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 166.640 586.335 167.240 ;
    END
  END pcpi_rs2[5]
  PIN pcpi_rs2[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 326.440 4.000 327.040 ;
    END
  END pcpi_rs2[6]
  PIN pcpi_rs2[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 13.640 586.335 14.240 ;
    END
  END pcpi_rs2[7]
  PIN pcpi_rs2[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 93.470 0.000 93.750 4.000 ;
    END
  END pcpi_rs2[8]
  PIN pcpi_rs2[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 286.670 0.000 286.950 4.000 ;
    END
  END pcpi_rs2[9]
  PIN pcpi_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 251.640 586.335 252.240 ;
    END
  END pcpi_valid
  PIN pcpi_wait
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 466.990 593.055 467.270 597.055 ;
    END
  END pcpi_wait
  PIN pcpi_wr
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 530.440 586.335 531.040 ;
    END
  END pcpi_wr
  PIN resetn
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 17.040 586.335 17.640 ;
    END
  END resetn
  PIN trace_data[0]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 45.170 0.000 45.450 4.000 ;
    END
  END trace_data[0]
  PIN trace_data[10]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 333.240 586.335 333.840 ;
    END
  END trace_data[10]
  PIN trace_data[11]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 9.750 0.000 10.030 4.000 ;
    END
  END trace_data[11]
  PIN trace_data[12]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 547.440 586.335 548.040 ;
    END
  END trace_data[12]
  PIN trace_data[13]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 444.450 593.055 444.730 597.055 ;
    END
  END trace_data[13]
  PIN trace_data[14]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 61.240 586.335 61.840 ;
    END
  END trace_data[14]
  PIN trace_data[15]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 425.130 593.055 425.410 597.055 ;
    END
  END trace_data[15]
  PIN trace_data[16]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 170.040 4.000 170.640 ;
    END
  END trace_data[16]
  PIN trace_data[17]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 190.440 4.000 191.040 ;
    END
  END trace_data[17]
  PIN trace_data[18]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 389.710 0.000 389.990 4.000 ;
    END
  END trace_data[18]
  PIN trace_data[19]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 0.090 0.000 0.370 4.000 ;
    END
  END trace_data[19]
  PIN trace_data[1]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 457.330 0.000 457.610 4.000 ;
    END
  END trace_data[1]
  PIN trace_data[20]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 289.040 4.000 289.640 ;
    END
  END trace_data[20]
  PIN trace_data[21]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 530.440 4.000 531.040 ;
    END
  END trace_data[21]
  PIN trace_data[22]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 170.750 593.055 171.030 597.055 ;
    END
  END trace_data[22]
  PIN trace_data[23]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 200.640 4.000 201.240 ;
    END
  END trace_data[23]
  PIN trace_data[24]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 116.010 0.000 116.290 4.000 ;
    END
  END trace_data[24]
  PIN trace_data[25]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 38.730 0.000 39.010 4.000 ;
    END
  END trace_data[25]
  PIN trace_data[26]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 593.055 309.490 597.055 ;
    END
  END trace_data[26]
  PIN trace_data[27]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 177.190 593.055 177.470 597.055 ;
    END
  END trace_data[27]
  PIN trace_data[28]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 309.210 0.000 309.490 4.000 ;
    END
  END trace_data[28]
  PIN trace_data[29]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 409.030 593.055 409.310 597.055 ;
    END
  END trace_data[29]
  PIN trace_data[2]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 159.840 586.335 160.440 ;
    END
  END trace_data[2]
  PIN trace_data[30]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 397.840 4.000 398.440 ;
    END
  END trace_data[30]
  PIN trace_data[31]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 459.040 586.335 459.640 ;
    END
  END trace_data[31]
  PIN trace_data[32]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 128.890 0.000 129.170 4.000 ;
    END
  END trace_data[32]
  PIN trace_data[33]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 219.050 0.000 219.330 4.000 ;
    END
  END trace_data[33]
  PIN trace_data[34]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 51.040 4.000 51.640 ;
    END
  END trace_data[34]
  PIN trace_data[35]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 435.240 586.335 435.840 ;
    END
  END trace_data[35]
  PIN trace_data[3]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 347.850 0.000 348.130 4.000 ;
    END
  END trace_data[3]
  PIN trace_data[4]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 386.490 593.055 386.770 597.055 ;
    END
  END trace_data[4]
  PIN trace_data[5]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 380.050 593.055 380.330 597.055 ;
    END
  END trace_data[5]
  PIN trace_data[6]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 557.640 4.000 558.240 ;
    END
  END trace_data[6]
  PIN trace_data[7]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 70.930 593.055 71.210 597.055 ;
    END
  END trace_data[7]
  PIN trace_data[8]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT 415.470 0.000 415.750 4.000 ;
    END
  END trace_data[8]
  PIN trace_data[9]
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 136.040 4.000 136.640 ;
    END
  END trace_data[9]
  PIN trace_valid
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 0.000 499.840 4.000 500.440 ;
    END
  END trace_valid
  PIN trap
    DIRECTION OUTPUT TRISTATE ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT 582.335 285.640 586.335 286.240 ;
    END
  END trap
  OBS
      LAYER li1 ;
        RECT 5.520 10.795 580.520 584.885 ;
      LAYER met1 ;
        RECT 0.070 277.340 586.335 593.600 ;
        RECT 0.070 275.840 586.340 277.340 ;
        RECT 0.070 5.820 586.335 275.840 ;
      LAYER met2 ;
        RECT 0.100 592.775 3.030 595.525 ;
        RECT 3.870 592.775 6.250 595.525 ;
        RECT 7.090 592.775 12.690 595.525 ;
        RECT 13.530 592.775 19.130 595.525 ;
        RECT 19.970 592.775 25.570 595.525 ;
        RECT 26.410 592.775 32.010 595.525 ;
        RECT 32.850 592.775 35.230 595.525 ;
        RECT 36.070 592.775 41.670 595.525 ;
        RECT 42.510 592.775 48.110 595.525 ;
        RECT 48.950 592.775 54.550 595.525 ;
        RECT 55.390 592.775 57.770 595.525 ;
        RECT 58.610 592.775 64.210 595.525 ;
        RECT 65.050 592.775 70.650 595.525 ;
        RECT 71.490 592.775 77.090 595.525 ;
        RECT 77.930 592.775 80.310 595.525 ;
        RECT 81.150 592.775 86.750 595.525 ;
        RECT 87.590 592.775 93.190 595.525 ;
        RECT 94.030 592.775 99.630 595.525 ;
        RECT 100.470 592.775 102.850 595.525 ;
        RECT 103.690 592.775 109.290 595.525 ;
        RECT 110.130 592.775 115.730 595.525 ;
        RECT 116.570 592.775 122.170 595.525 ;
        RECT 123.010 592.775 125.390 595.525 ;
        RECT 126.230 592.775 131.830 595.525 ;
        RECT 132.670 592.775 138.270 595.525 ;
        RECT 139.110 592.775 144.710 595.525 ;
        RECT 145.550 592.775 147.930 595.525 ;
        RECT 148.770 592.775 154.370 595.525 ;
        RECT 155.210 592.775 160.810 595.525 ;
        RECT 161.650 592.775 167.250 595.525 ;
        RECT 168.090 592.775 170.470 595.525 ;
        RECT 171.310 592.775 176.910 595.525 ;
        RECT 177.750 592.775 183.350 595.525 ;
        RECT 184.190 592.775 189.790 595.525 ;
        RECT 190.630 592.775 193.010 595.525 ;
        RECT 193.850 592.775 199.450 595.525 ;
        RECT 200.290 592.775 205.890 595.525 ;
        RECT 206.730 592.775 212.330 595.525 ;
        RECT 213.170 592.775 215.550 595.525 ;
        RECT 216.390 592.775 221.990 595.525 ;
        RECT 222.830 592.775 228.430 595.525 ;
        RECT 229.270 592.775 234.870 595.525 ;
        RECT 235.710 592.775 238.090 595.525 ;
        RECT 238.930 592.775 244.530 595.525 ;
        RECT 245.370 592.775 250.970 595.525 ;
        RECT 251.810 592.775 257.410 595.525 ;
        RECT 258.250 592.775 260.630 595.525 ;
        RECT 261.470 592.775 267.070 595.525 ;
        RECT 267.910 592.775 273.510 595.525 ;
        RECT 274.350 592.775 279.950 595.525 ;
        RECT 280.790 592.775 283.170 595.525 ;
        RECT 284.010 592.775 289.610 595.525 ;
        RECT 290.450 592.775 296.050 595.525 ;
        RECT 296.890 592.775 302.490 595.525 ;
        RECT 303.330 592.775 308.930 595.525 ;
        RECT 309.770 592.775 312.150 595.525 ;
        RECT 312.990 592.775 318.590 595.525 ;
        RECT 319.430 592.775 325.030 595.525 ;
        RECT 325.870 592.775 331.470 595.525 ;
        RECT 332.310 592.775 334.690 595.525 ;
        RECT 335.530 592.775 341.130 595.525 ;
        RECT 341.970 592.775 347.570 595.525 ;
        RECT 348.410 592.775 354.010 595.525 ;
        RECT 354.850 592.775 357.230 595.525 ;
        RECT 358.070 592.775 363.670 595.525 ;
        RECT 364.510 592.775 370.110 595.525 ;
        RECT 370.950 592.775 376.550 595.525 ;
        RECT 377.390 592.775 379.770 595.525 ;
        RECT 380.610 592.775 386.210 595.525 ;
        RECT 387.050 592.775 392.650 595.525 ;
        RECT 393.490 592.775 399.090 595.525 ;
        RECT 399.930 592.775 402.310 595.525 ;
        RECT 403.150 592.775 408.750 595.525 ;
        RECT 409.590 592.775 415.190 595.525 ;
        RECT 416.030 592.775 421.630 595.525 ;
        RECT 422.470 592.775 424.850 595.525 ;
        RECT 425.690 592.775 431.290 595.525 ;
        RECT 432.130 592.775 437.730 595.525 ;
        RECT 438.570 592.775 444.170 595.525 ;
        RECT 445.010 592.775 447.390 595.525 ;
        RECT 448.230 592.775 453.830 595.525 ;
        RECT 454.670 592.775 460.270 595.525 ;
        RECT 461.110 592.775 466.710 595.525 ;
        RECT 467.550 592.775 469.930 595.525 ;
        RECT 470.770 592.775 476.370 595.525 ;
        RECT 477.210 592.775 482.810 595.525 ;
        RECT 483.650 592.775 489.250 595.525 ;
        RECT 490.090 592.775 492.470 595.525 ;
        RECT 493.310 592.775 498.910 595.525 ;
        RECT 499.750 592.775 505.350 595.525 ;
        RECT 506.190 592.775 511.790 595.525 ;
        RECT 512.630 592.775 515.010 595.525 ;
        RECT 515.850 592.775 521.450 595.525 ;
        RECT 522.290 592.775 527.890 595.525 ;
        RECT 528.730 592.775 534.330 595.525 ;
        RECT 535.170 592.775 537.550 595.525 ;
        RECT 538.390 592.775 543.990 595.525 ;
        RECT 544.830 592.775 550.430 595.525 ;
        RECT 551.270 592.775 556.870 595.525 ;
        RECT 557.710 592.775 560.090 595.525 ;
        RECT 560.930 592.775 566.530 595.525 ;
        RECT 567.370 592.775 572.970 595.525 ;
        RECT 573.810 592.775 579.410 595.525 ;
        RECT 580.250 592.775 582.630 595.525 ;
        RECT 583.470 592.775 586.335 595.525 ;
        RECT 0.100 496.870 586.335 592.775 ;
        RECT 0.100 393.820 586.340 496.870 ;
        RECT 0.100 338.170 586.335 393.820 ;
        RECT 0.100 276.520 586.340 338.170 ;
        RECT 0.100 4.280 586.335 276.520 ;
        RECT 0.650 0.155 3.030 4.280 ;
        RECT 3.870 0.155 9.470 4.280 ;
        RECT 10.310 0.155 15.910 4.280 ;
        RECT 16.750 0.155 22.350 4.280 ;
        RECT 23.190 0.155 25.570 4.280 ;
        RECT 26.410 0.155 32.010 4.280 ;
        RECT 32.850 0.155 38.450 4.280 ;
        RECT 39.290 0.155 44.890 4.280 ;
        RECT 45.730 0.155 48.110 4.280 ;
        RECT 48.950 0.155 54.550 4.280 ;
        RECT 55.390 0.155 60.990 4.280 ;
        RECT 61.830 0.155 67.430 4.280 ;
        RECT 68.270 0.155 70.650 4.280 ;
        RECT 71.490 0.155 77.090 4.280 ;
        RECT 77.930 0.155 83.530 4.280 ;
        RECT 84.370 0.155 89.970 4.280 ;
        RECT 90.810 0.155 93.190 4.280 ;
        RECT 94.030 0.155 99.630 4.280 ;
        RECT 100.470 0.155 106.070 4.280 ;
        RECT 106.910 0.155 112.510 4.280 ;
        RECT 113.350 0.155 115.730 4.280 ;
        RECT 116.570 0.155 122.170 4.280 ;
        RECT 123.010 0.155 128.610 4.280 ;
        RECT 129.450 0.155 135.050 4.280 ;
        RECT 135.890 0.155 138.270 4.280 ;
        RECT 139.110 0.155 144.710 4.280 ;
        RECT 145.550 0.155 151.150 4.280 ;
        RECT 151.990 0.155 157.590 4.280 ;
        RECT 158.430 0.155 160.810 4.280 ;
        RECT 161.650 0.155 167.250 4.280 ;
        RECT 168.090 0.155 173.690 4.280 ;
        RECT 174.530 0.155 180.130 4.280 ;
        RECT 180.970 0.155 183.350 4.280 ;
        RECT 184.190 0.155 189.790 4.280 ;
        RECT 190.630 0.155 196.230 4.280 ;
        RECT 197.070 0.155 202.670 4.280 ;
        RECT 203.510 0.155 205.890 4.280 ;
        RECT 206.730 0.155 212.330 4.280 ;
        RECT 213.170 0.155 218.770 4.280 ;
        RECT 219.610 0.155 225.210 4.280 ;
        RECT 226.050 0.155 228.430 4.280 ;
        RECT 229.270 0.155 234.870 4.280 ;
        RECT 235.710 0.155 241.310 4.280 ;
        RECT 242.150 0.155 247.750 4.280 ;
        RECT 248.590 0.155 250.970 4.280 ;
        RECT 251.810 0.155 257.410 4.280 ;
        RECT 258.250 0.155 263.850 4.280 ;
        RECT 264.690 0.155 270.290 4.280 ;
        RECT 271.130 0.155 273.510 4.280 ;
        RECT 274.350 0.155 279.950 4.280 ;
        RECT 280.790 0.155 286.390 4.280 ;
        RECT 287.230 0.155 292.830 4.280 ;
        RECT 293.670 0.155 299.270 4.280 ;
        RECT 300.110 0.155 302.490 4.280 ;
        RECT 303.330 0.155 308.930 4.280 ;
        RECT 309.770 0.155 315.370 4.280 ;
        RECT 316.210 0.155 321.810 4.280 ;
        RECT 322.650 0.155 325.030 4.280 ;
        RECT 325.870 0.155 331.470 4.280 ;
        RECT 332.310 0.155 337.910 4.280 ;
        RECT 338.750 0.155 344.350 4.280 ;
        RECT 345.190 0.155 347.570 4.280 ;
        RECT 348.410 0.155 354.010 4.280 ;
        RECT 354.850 0.155 360.450 4.280 ;
        RECT 361.290 0.155 366.890 4.280 ;
        RECT 367.730 0.155 370.110 4.280 ;
        RECT 370.950 0.155 376.550 4.280 ;
        RECT 377.390 0.155 382.990 4.280 ;
        RECT 383.830 0.155 389.430 4.280 ;
        RECT 390.270 0.155 392.650 4.280 ;
        RECT 393.490 0.155 399.090 4.280 ;
        RECT 399.930 0.155 405.530 4.280 ;
        RECT 406.370 0.155 411.970 4.280 ;
        RECT 412.810 0.155 415.190 4.280 ;
        RECT 416.030 0.155 421.630 4.280 ;
        RECT 422.470 0.155 428.070 4.280 ;
        RECT 428.910 0.155 434.510 4.280 ;
        RECT 435.350 0.155 437.730 4.280 ;
        RECT 438.570 0.155 444.170 4.280 ;
        RECT 445.010 0.155 450.610 4.280 ;
        RECT 451.450 0.155 457.050 4.280 ;
        RECT 457.890 0.155 460.270 4.280 ;
        RECT 461.110 0.155 466.710 4.280 ;
        RECT 467.550 0.155 473.150 4.280 ;
        RECT 473.990 0.155 479.590 4.280 ;
        RECT 480.430 0.155 482.810 4.280 ;
        RECT 483.650 0.155 489.250 4.280 ;
        RECT 490.090 0.155 495.690 4.280 ;
        RECT 496.530 0.155 502.130 4.280 ;
        RECT 502.970 0.155 505.350 4.280 ;
        RECT 506.190 0.155 511.790 4.280 ;
        RECT 512.630 0.155 518.230 4.280 ;
        RECT 519.070 0.155 524.670 4.280 ;
        RECT 525.510 0.155 527.890 4.280 ;
        RECT 528.730 0.155 534.330 4.280 ;
        RECT 535.170 0.155 540.770 4.280 ;
        RECT 541.610 0.155 547.210 4.280 ;
        RECT 548.050 0.155 550.430 4.280 ;
        RECT 551.270 0.155 556.870 4.280 ;
        RECT 557.710 0.155 563.310 4.280 ;
        RECT 564.150 0.155 569.750 4.280 ;
        RECT 570.590 0.155 576.190 4.280 ;
        RECT 577.030 0.155 579.410 4.280 ;
        RECT 580.250 0.155 586.335 4.280 ;
      LAYER met3 ;
        RECT 4.400 594.640 585.975 595.505 ;
        RECT 2.825 592.640 585.975 594.640 ;
        RECT 2.825 591.240 581.935 592.640 ;
        RECT 2.825 589.240 585.975 591.240 ;
        RECT 4.400 587.840 585.975 589.240 ;
        RECT 2.825 585.840 585.975 587.840 ;
        RECT 2.825 584.440 581.935 585.840 ;
        RECT 2.825 582.440 585.975 584.440 ;
        RECT 4.400 581.040 585.975 582.440 ;
        RECT 2.825 579.040 585.975 581.040 ;
        RECT 4.400 577.640 581.935 579.040 ;
        RECT 2.825 572.240 585.975 577.640 ;
        RECT 4.400 570.840 581.935 572.240 ;
        RECT 2.825 568.840 585.975 570.840 ;
        RECT 2.825 567.440 581.935 568.840 ;
        RECT 2.825 565.440 585.975 567.440 ;
        RECT 4.400 564.040 585.975 565.440 ;
        RECT 2.825 562.040 585.975 564.040 ;
        RECT 2.825 560.640 581.935 562.040 ;
        RECT 2.825 558.640 585.975 560.640 ;
        RECT 4.400 557.240 585.975 558.640 ;
        RECT 2.825 555.240 585.975 557.240 ;
        RECT 4.400 553.840 581.935 555.240 ;
        RECT 2.825 548.440 585.975 553.840 ;
        RECT 4.400 547.040 581.935 548.440 ;
        RECT 2.825 545.040 585.975 547.040 ;
        RECT 2.825 543.640 581.935 545.040 ;
        RECT 2.825 541.640 585.975 543.640 ;
        RECT 4.400 540.240 585.975 541.640 ;
        RECT 2.825 538.240 585.975 540.240 ;
        RECT 2.825 536.840 581.935 538.240 ;
        RECT 2.825 534.840 585.975 536.840 ;
        RECT 4.400 533.440 585.975 534.840 ;
        RECT 2.825 531.440 585.975 533.440 ;
        RECT 4.400 530.040 581.935 531.440 ;
        RECT 2.825 524.640 585.975 530.040 ;
        RECT 4.400 523.240 581.935 524.640 ;
        RECT 2.825 521.240 585.975 523.240 ;
        RECT 2.825 519.840 581.935 521.240 ;
        RECT 2.825 517.840 585.975 519.840 ;
        RECT 4.400 516.440 585.975 517.840 ;
        RECT 2.825 514.440 585.975 516.440 ;
        RECT 2.825 513.040 581.935 514.440 ;
        RECT 2.825 511.040 585.975 513.040 ;
        RECT 4.400 509.640 585.975 511.040 ;
        RECT 2.825 507.640 585.975 509.640 ;
        RECT 4.400 506.240 581.935 507.640 ;
        RECT 2.825 500.840 585.975 506.240 ;
        RECT 4.400 499.440 581.935 500.840 ;
        RECT 2.825 497.440 585.975 499.440 ;
        RECT 2.825 496.040 581.935 497.440 ;
        RECT 2.825 494.040 585.975 496.040 ;
        RECT 4.400 492.640 585.975 494.040 ;
        RECT 2.825 490.640 585.975 492.640 ;
        RECT 2.825 489.240 581.935 490.640 ;
        RECT 2.825 487.240 585.975 489.240 ;
        RECT 4.400 485.840 585.975 487.240 ;
        RECT 2.825 483.840 585.975 485.840 ;
        RECT 4.400 482.440 581.935 483.840 ;
        RECT 2.825 477.040 585.975 482.440 ;
        RECT 4.400 475.640 581.935 477.040 ;
        RECT 2.825 473.640 585.975 475.640 ;
        RECT 2.825 472.240 581.935 473.640 ;
        RECT 2.825 470.240 585.975 472.240 ;
        RECT 4.400 468.840 585.975 470.240 ;
        RECT 2.825 466.840 585.975 468.840 ;
        RECT 2.825 465.440 581.935 466.840 ;
        RECT 2.825 463.440 585.975 465.440 ;
        RECT 4.400 462.040 585.975 463.440 ;
        RECT 2.825 460.040 585.975 462.040 ;
        RECT 4.400 458.640 581.935 460.040 ;
        RECT 2.825 453.240 585.975 458.640 ;
        RECT 4.400 451.840 581.935 453.240 ;
        RECT 2.825 449.840 585.975 451.840 ;
        RECT 2.825 448.440 581.935 449.840 ;
        RECT 2.825 446.440 585.975 448.440 ;
        RECT 4.400 445.040 585.975 446.440 ;
        RECT 2.825 443.040 585.975 445.040 ;
        RECT 2.825 441.640 581.935 443.040 ;
        RECT 2.825 439.640 585.975 441.640 ;
        RECT 4.400 438.240 585.975 439.640 ;
        RECT 2.825 436.240 585.975 438.240 ;
        RECT 4.400 434.840 581.935 436.240 ;
        RECT 2.825 429.440 585.975 434.840 ;
        RECT 4.400 428.040 581.935 429.440 ;
        RECT 2.825 426.040 585.975 428.040 ;
        RECT 2.825 424.640 581.935 426.040 ;
        RECT 2.825 422.640 585.975 424.640 ;
        RECT 4.400 421.240 585.975 422.640 ;
        RECT 2.825 419.240 585.975 421.240 ;
        RECT 2.825 417.840 581.935 419.240 ;
        RECT 2.825 415.840 585.975 417.840 ;
        RECT 4.400 414.440 585.975 415.840 ;
        RECT 2.825 412.440 585.975 414.440 ;
        RECT 4.400 411.040 581.935 412.440 ;
        RECT 2.825 405.640 585.975 411.040 ;
        RECT 4.400 404.240 581.935 405.640 ;
        RECT 2.825 402.240 585.975 404.240 ;
        RECT 2.825 400.840 581.935 402.240 ;
        RECT 2.825 398.840 585.975 400.840 ;
        RECT 4.400 397.440 585.975 398.840 ;
        RECT 2.825 395.440 585.975 397.440 ;
        RECT 2.825 394.040 581.935 395.440 ;
        RECT 2.825 392.040 585.975 394.040 ;
        RECT 4.400 390.640 585.975 392.040 ;
        RECT 2.825 388.640 585.975 390.640 ;
        RECT 4.400 387.240 581.935 388.640 ;
        RECT 2.825 381.840 585.975 387.240 ;
        RECT 4.400 380.440 581.935 381.840 ;
        RECT 2.825 378.440 585.975 380.440 ;
        RECT 2.825 377.040 581.935 378.440 ;
        RECT 2.825 375.040 585.975 377.040 ;
        RECT 4.400 373.640 585.975 375.040 ;
        RECT 2.825 371.640 585.975 373.640 ;
        RECT 2.825 370.240 581.935 371.640 ;
        RECT 2.825 368.240 585.975 370.240 ;
        RECT 4.400 366.840 585.975 368.240 ;
        RECT 2.825 364.840 585.975 366.840 ;
        RECT 4.400 363.440 581.935 364.840 ;
        RECT 2.825 358.040 585.975 363.440 ;
        RECT 4.400 356.640 581.935 358.040 ;
        RECT 2.825 354.640 585.975 356.640 ;
        RECT 2.825 353.240 581.935 354.640 ;
        RECT 2.825 351.240 585.975 353.240 ;
        RECT 4.400 349.840 585.975 351.240 ;
        RECT 2.825 347.840 585.975 349.840 ;
        RECT 2.825 346.440 581.935 347.840 ;
        RECT 2.825 344.440 585.975 346.440 ;
        RECT 4.400 343.040 585.975 344.440 ;
        RECT 2.825 341.040 585.975 343.040 ;
        RECT 4.400 339.640 581.935 341.040 ;
        RECT 2.825 334.240 585.975 339.640 ;
        RECT 4.400 332.840 581.935 334.240 ;
        RECT 2.825 330.840 585.975 332.840 ;
        RECT 2.825 329.440 581.935 330.840 ;
        RECT 2.825 327.440 585.975 329.440 ;
        RECT 4.400 326.040 585.975 327.440 ;
        RECT 2.825 324.040 585.975 326.040 ;
        RECT 2.825 322.640 581.935 324.040 ;
        RECT 2.825 320.640 585.975 322.640 ;
        RECT 4.400 319.240 585.975 320.640 ;
        RECT 2.825 317.240 585.975 319.240 ;
        RECT 4.400 315.840 581.935 317.240 ;
        RECT 2.825 310.440 585.975 315.840 ;
        RECT 4.400 309.040 581.935 310.440 ;
        RECT 2.825 307.040 585.975 309.040 ;
        RECT 2.825 305.640 581.935 307.040 ;
        RECT 2.825 303.640 585.975 305.640 ;
        RECT 4.400 302.240 585.975 303.640 ;
        RECT 2.825 300.240 585.975 302.240 ;
        RECT 2.825 298.840 581.935 300.240 ;
        RECT 2.825 296.840 585.975 298.840 ;
        RECT 4.400 295.440 585.975 296.840 ;
        RECT 2.825 293.440 585.975 295.440 ;
        RECT 2.825 292.040 581.935 293.440 ;
        RECT 2.825 290.040 585.975 292.040 ;
        RECT 4.400 288.640 585.975 290.040 ;
        RECT 2.825 286.640 585.975 288.640 ;
        RECT 4.400 285.240 581.935 286.640 ;
        RECT 2.825 279.840 585.975 285.240 ;
        RECT 4.400 278.440 581.935 279.840 ;
        RECT 2.825 276.440 585.975 278.440 ;
        RECT 2.825 275.040 581.935 276.440 ;
        RECT 2.825 273.040 585.975 275.040 ;
        RECT 4.400 271.640 585.975 273.040 ;
        RECT 2.825 269.640 585.975 271.640 ;
        RECT 2.825 268.240 581.935 269.640 ;
        RECT 2.825 266.240 585.975 268.240 ;
        RECT 4.400 264.840 585.975 266.240 ;
        RECT 2.825 262.840 585.975 264.840 ;
        RECT 4.400 261.440 581.935 262.840 ;
        RECT 2.825 256.040 585.975 261.440 ;
        RECT 4.400 254.640 581.935 256.040 ;
        RECT 2.825 252.640 585.975 254.640 ;
        RECT 2.825 251.240 581.935 252.640 ;
        RECT 2.825 249.240 585.975 251.240 ;
        RECT 4.400 247.840 585.975 249.240 ;
        RECT 2.825 245.840 585.975 247.840 ;
        RECT 2.825 244.440 581.935 245.840 ;
        RECT 2.825 242.440 585.975 244.440 ;
        RECT 4.400 241.040 585.975 242.440 ;
        RECT 2.825 239.040 585.975 241.040 ;
        RECT 4.400 237.640 581.935 239.040 ;
        RECT 2.825 232.240 585.975 237.640 ;
        RECT 4.400 230.840 581.935 232.240 ;
        RECT 2.825 228.840 585.975 230.840 ;
        RECT 2.825 227.440 581.935 228.840 ;
        RECT 2.825 225.440 585.975 227.440 ;
        RECT 4.400 224.040 585.975 225.440 ;
        RECT 2.825 222.040 585.975 224.040 ;
        RECT 2.825 220.640 581.935 222.040 ;
        RECT 2.825 218.640 585.975 220.640 ;
        RECT 4.400 217.240 585.975 218.640 ;
        RECT 2.825 215.240 585.975 217.240 ;
        RECT 4.400 213.840 581.935 215.240 ;
        RECT 2.825 208.440 585.975 213.840 ;
        RECT 4.400 207.040 581.935 208.440 ;
        RECT 2.825 205.040 585.975 207.040 ;
        RECT 2.825 203.640 581.935 205.040 ;
        RECT 2.825 201.640 585.975 203.640 ;
        RECT 4.400 200.240 585.975 201.640 ;
        RECT 2.825 198.240 585.975 200.240 ;
        RECT 2.825 196.840 581.935 198.240 ;
        RECT 2.825 194.840 585.975 196.840 ;
        RECT 4.400 193.440 585.975 194.840 ;
        RECT 2.825 191.440 585.975 193.440 ;
        RECT 4.400 190.040 581.935 191.440 ;
        RECT 2.825 184.640 585.975 190.040 ;
        RECT 4.400 183.240 581.935 184.640 ;
        RECT 2.825 181.240 585.975 183.240 ;
        RECT 2.825 179.840 581.935 181.240 ;
        RECT 2.825 177.840 585.975 179.840 ;
        RECT 4.400 176.440 585.975 177.840 ;
        RECT 2.825 174.440 585.975 176.440 ;
        RECT 2.825 173.040 581.935 174.440 ;
        RECT 2.825 171.040 585.975 173.040 ;
        RECT 4.400 169.640 585.975 171.040 ;
        RECT 2.825 167.640 585.975 169.640 ;
        RECT 4.400 166.240 581.935 167.640 ;
        RECT 2.825 160.840 585.975 166.240 ;
        RECT 4.400 159.440 581.935 160.840 ;
        RECT 2.825 157.440 585.975 159.440 ;
        RECT 2.825 156.040 581.935 157.440 ;
        RECT 2.825 154.040 585.975 156.040 ;
        RECT 4.400 152.640 585.975 154.040 ;
        RECT 2.825 150.640 585.975 152.640 ;
        RECT 2.825 149.240 581.935 150.640 ;
        RECT 2.825 147.240 585.975 149.240 ;
        RECT 4.400 145.840 585.975 147.240 ;
        RECT 2.825 143.840 585.975 145.840 ;
        RECT 4.400 142.440 581.935 143.840 ;
        RECT 2.825 137.040 585.975 142.440 ;
        RECT 4.400 135.640 581.935 137.040 ;
        RECT 2.825 133.640 585.975 135.640 ;
        RECT 2.825 132.240 581.935 133.640 ;
        RECT 2.825 130.240 585.975 132.240 ;
        RECT 4.400 128.840 585.975 130.240 ;
        RECT 2.825 126.840 585.975 128.840 ;
        RECT 2.825 125.440 581.935 126.840 ;
        RECT 2.825 123.440 585.975 125.440 ;
        RECT 4.400 122.040 585.975 123.440 ;
        RECT 2.825 120.040 585.975 122.040 ;
        RECT 4.400 118.640 581.935 120.040 ;
        RECT 2.825 113.240 585.975 118.640 ;
        RECT 4.400 111.840 581.935 113.240 ;
        RECT 2.825 109.840 585.975 111.840 ;
        RECT 2.825 108.440 581.935 109.840 ;
        RECT 2.825 106.440 585.975 108.440 ;
        RECT 4.400 105.040 585.975 106.440 ;
        RECT 2.825 103.040 585.975 105.040 ;
        RECT 2.825 101.640 581.935 103.040 ;
        RECT 2.825 99.640 585.975 101.640 ;
        RECT 4.400 98.240 585.975 99.640 ;
        RECT 2.825 96.240 585.975 98.240 ;
        RECT 4.400 94.840 581.935 96.240 ;
        RECT 2.825 89.440 585.975 94.840 ;
        RECT 4.400 88.040 581.935 89.440 ;
        RECT 2.825 86.040 585.975 88.040 ;
        RECT 2.825 84.640 581.935 86.040 ;
        RECT 2.825 82.640 585.975 84.640 ;
        RECT 4.400 81.240 585.975 82.640 ;
        RECT 2.825 79.240 585.975 81.240 ;
        RECT 2.825 77.840 581.935 79.240 ;
        RECT 2.825 75.840 585.975 77.840 ;
        RECT 4.400 74.440 585.975 75.840 ;
        RECT 2.825 72.440 585.975 74.440 ;
        RECT 4.400 71.040 581.935 72.440 ;
        RECT 2.825 65.640 585.975 71.040 ;
        RECT 4.400 64.240 581.935 65.640 ;
        RECT 2.825 62.240 585.975 64.240 ;
        RECT 2.825 60.840 581.935 62.240 ;
        RECT 2.825 58.840 585.975 60.840 ;
        RECT 4.400 57.440 585.975 58.840 ;
        RECT 2.825 55.440 585.975 57.440 ;
        RECT 2.825 54.040 581.935 55.440 ;
        RECT 2.825 52.040 585.975 54.040 ;
        RECT 4.400 50.640 585.975 52.040 ;
        RECT 2.825 48.640 585.975 50.640 ;
        RECT 4.400 47.240 581.935 48.640 ;
        RECT 2.825 41.840 585.975 47.240 ;
        RECT 4.400 40.440 581.935 41.840 ;
        RECT 2.825 38.440 585.975 40.440 ;
        RECT 2.825 37.040 581.935 38.440 ;
        RECT 2.825 35.040 585.975 37.040 ;
        RECT 4.400 33.640 585.975 35.040 ;
        RECT 2.825 31.640 585.975 33.640 ;
        RECT 2.825 30.240 581.935 31.640 ;
        RECT 2.825 28.240 585.975 30.240 ;
        RECT 4.400 26.840 585.975 28.240 ;
        RECT 2.825 24.840 585.975 26.840 ;
        RECT 4.400 23.440 581.935 24.840 ;
        RECT 2.825 18.040 585.975 23.440 ;
        RECT 4.400 16.640 581.935 18.040 ;
        RECT 2.825 14.640 585.975 16.640 ;
        RECT 2.825 13.240 581.935 14.640 ;
        RECT 2.825 11.240 585.975 13.240 ;
        RECT 4.400 9.840 585.975 11.240 ;
        RECT 2.825 7.840 585.975 9.840 ;
        RECT 2.825 6.440 581.935 7.840 ;
        RECT 2.825 4.440 585.975 6.440 ;
        RECT 4.400 3.040 585.975 4.440 ;
        RECT 2.825 1.040 585.975 3.040 ;
        RECT 2.825 0.175 581.935 1.040 ;
      LAYER met4 ;
        RECT 7.655 12.415 20.640 584.625 ;
        RECT 23.040 12.415 97.440 584.625 ;
        RECT 99.840 12.415 174.240 584.625 ;
        RECT 176.640 12.415 251.040 584.625 ;
        RECT 253.440 12.415 327.840 584.625 ;
        RECT 330.240 12.415 404.640 584.625 ;
        RECT 407.040 12.415 481.440 584.625 ;
        RECT 483.840 12.415 558.240 584.625 ;
        RECT 560.640 12.415 582.065 584.625 ;
      LAYER met5 ;
        RECT 36.460 565.820 574.420 570.300 ;
        RECT 36.460 489.230 574.420 561.020 ;
        RECT 36.460 412.640 574.420 484.430 ;
        RECT 36.460 336.050 574.420 407.840 ;
        RECT 36.460 259.460 574.420 331.250 ;
        RECT 36.460 182.870 574.420 254.660 ;
        RECT 36.460 106.300 574.420 178.070 ;
  END
END picorv32_woready
END LIBRARY

